package AES_Package;
import uvm_pkg::*;
parameter Encrypt_count =100;
 `include"uvm_macros.svh"
 `include "AES_seq_item.sv"
 `include "AES_Sequancer.sv"
 `include "AES_Driver.sv"   
 `include "AES_Monitor.sv"
 `include "AES_Agent.sv"
 `include "AES_Scoreboard.sv"
 `include "AES_coverage_collector.sv"
 `include "AES_Sequance.sv"
 `include "AES_ENV.sv"
 `include "AES_TEST.sv"
endpackage
