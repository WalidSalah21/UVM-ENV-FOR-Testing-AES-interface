interface  AES_INTERFACE();
    logic [127:0]  in ;
    logic [127:0]  key;
    logic [127:0]  out;
endinterface
